LIBRARY ieee;
USE ieee.std_logic_1164.all;
ENTITY HDU IS
GENERIC (n : integer := 3); 
PORT(Is_Load, Has_SRC2,Has_SRC1:IN STD_LOGIC;
SRC2_ADD,SRC1_ADD,LDD_ADD:IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
Is_Hazard: OUT STD_LOGIC);     
END HDU;

ARCHITECTURE MY_HDU OF HDU IS
  BEGIN
Is_Hazard <= '1' WHEN Is_Load = '1' AND Has_SRC2 = '1' AND LDD_ADD = SRC2_ADD
ELSE '1' WHEN Is_Load = '1' AND Has_SRC1 = '1' AND LDD_ADD = SRC1_ADD
ELSE '0'; 
  
END ARCHITECTURE;